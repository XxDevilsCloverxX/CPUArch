`timescale 1ns / 1ps

/*
Name: Silas Rodriguez
R-Number: R-11679913
Assignment: Project 6
*/

/**

    * DataPath.v
    * This module is responsible for organizing the CPU architecthure and connecting all the modules together.
    
    * Inputs:
    *  clk - External Clock signal
    *  reset - External Reset signal
    
    * Outputs:
    *  None
*/
module CPU(
    input clk,      //clock
    input reset,    //reset
    output wire [31:0] GPR0, //General Purpose Register 0
);

    //create an instruction memory

    //create a program counter

    //create a register file

    //create an ALU

    //create a decoder

endmodule